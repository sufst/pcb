.title KiCad schematic
.model __NT6 
.model __J16 
.model __J14 
.model __J17 
.model __J13 
.model __J15 
.model __J11 
.model __SW2 
.model __NT3 
.model __NT4 
.model __SW1 
.model __J4 
.model __NT1 
.model __NT2 
.model __LV_GND1 
.model __J9 
.model __J10 
.model __J7 
.model __J5 
.model __J6 
.model __SW3 
.model __J8 
.model __NT5 
.model __J12 
.model __J3 
.model __J2 
.model __J1 
.model __J18 
.model __J19 
.model __J26 
.model __J30 
.model __J34 
.model __J29 
.model __J37 
.model __J35 
.model __J25 
.model __J24 
.model __J33 
.model __J32 
.model __J28 
.model __J31 
.model __J27 
.model __NT8 
.model __NT10 
.model __NT9 
.model __J36 
.model __J20 
.model __NT7 
.model __J22 
.model __J23 
.model __J21 
.model __J47 
.model __J46 
.model __J45 
.model __TSMP+.Resistor1 
.model __J38 
.model __TSMP-.Resistor1 
.model __J39 
.model __Discharge.Resistor1 
.model __J41 
.model __J40 
.model __J43 
.model __J44 
.model __J42 
.model __J48 
.model __J51 
.model __J49 
.model __J50 
.model __J54 
.model __J53 
.model __J52 
.model __J57 
.model __J56 
.model __J55 
.model __J58 
.model __J61 
.model __J60 
.model __J59 
.model __J66 
.model __J64 
.model __J65 
.model __J63 
.model __J62 
.model __TP2 
.model __TP1 
.model __J72 
.model __J76 
.model __J73 
.model __J77 
.model __J74 
.model __J78 
.model __J75 
.model __TP3 
.model __TP4 
.model __J70 
.model __J67 
.model __J71 
.model __J68 
.model __J69 
.model __SW4 
.model __D1 
.model __SW6 
.model __SW5 
.model __D4 
.model __D3 
.model __D2 
.model __J80 
.model __J79 
.model __J82 
.model __J81 
.model __BT1 
NT6 __NT6
J16 __J16
J14 __J14
J17 __J17
J13 __J13
J15 __J15
J11 __J11
SW2 __SW2
NT3 __NT3
NT4 __NT4
SW1 __SW1
J4 __J4
NT1 __NT1
NT2 __NT2
LV_GND1 __LV_GND1
J9 __J9
J10 __J10
J7 __J7
J5 __J5
J6 __J6
SW3 __SW3
J8 __J8
NT5 __NT5
J12 __J12
J3 __J3
J2 __J2
J1 __J1
J18 __J18
J19 __J19
J26 __J26
J30 __J30
J34 __J34
J29 __J29
J37 __J37
J35 __J35
J25 __J25
J24 __J24
J33 __J33
J32 __J32
J28 __J28
J31 __J31
J27 __J27
NT8 __NT8
NT10 __NT10
NT9 __NT9
J36 __J36
J20 __J20
NT7 __NT7
J22 __J22
J23 __J23
J21 __J21
J47 __J47
J46 __J46
J45 __J45
TSMP+.Resistor1 __TSMP+.Resistor1
J38 __J38
TSMP-.Resistor1 __TSMP-.Resistor1
J39 __J39
Discharge.Resistor1 __Discharge.Resistor1
J41 __J41
J40 __J40
J43 __J43
J44 __J44
J42 __J42
J48 __J48
J51 __J51
J49 __J49
J50 __J50
J54 __J54
J53 __J53
J52 __J52
J57 __J57
J56 __J56
J55 __J55
J58 __J58
J61 __J61
J60 __J60
J59 __J59
J66 __J66
J64 __J64
J65 __J65
J63 __J63
J62 __J62
TP2 __TP2
TP1 __TP1
R1 /Pedal Box/APPS.2.EXC /Pedal Box/APPS.1.EXC R_Small
J72 __J72
J76 __J76
J73 __J73
J77 __J77
J74 __J74
J78 __J78
J75 __J75
TP3 __TP3
TP4 __TP4
J70 __J70
J67 __J67
J71 __J71
J68 __J68
J69 __J69
SW4 __SW4
D1 __D1
SW6 __SW6
SW5 __SW5
D4 __D4
D3 __D3
D2 __D2
J80 __J80
J79 __J79
J82 __J82
J81 __J81
BT1 __BT1
.end
