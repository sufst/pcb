.title KiCad schematic
U2 Net-_D1-Pad2_ unconnected-_U2-Pad2_ unconnected-_U2-Pad3_ Net-_U1-Pad10_ unconnected-_U2-Pad5_ Net-_U1-Pad2_ Net-_U1-Pad4_ unconnected-_U2-Pad9_ Net-_U1-Pad10_ unconnected-_U2-Pad11_ unconnected-_U2-Pad12_ Net-_D2-Pad2_ 4013
U1 Net-_J1-Pad5_ Net-_U1-Pad2_ Net-_J1-Pad4_ Net-_U1-Pad4_ Net-_J1-Pad3_ Net-_U1-Pad6_ Net-_U1-Pad8_ Net-_J1-Pad2_ Net-_U1-Pad10_ /RESET 40106
U3 Net-_U1-Pad6_ unconnected-_U3-Pad9_ Net-_U1-Pad10_ unconnected-_U3-Pad11_ unconnected-_U3-Pad12_ Net-_D3-Pad2_ 4013
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ LED
R1 Net-_D1-Pad1_ GND R
U4 Net-_U1-Pad8_ unconnected-_U4-Pad9_ Net-_U1-Pad10_ unconnected-_U4-Pad11_ unconnected-_U4-Pad12_ Net-_D4-Pad2_ 4013
J1 /RESET Net-_J1-Pad2_ Net-_J1-Pad3_ Net-_J1-Pad4_ Net-_J1-Pad5_ Conn_01x05_Female
D2 Net-_D2-Pad1_ Net-_D2-Pad2_ LED
R2 Net-_D2-Pad1_ GND R
U5 /OUT Net-_D1-Pad2_ Net-_D2-Pad2_ Net-_D3-Pad2_ Net-_D4-Pad2_ 4072
R5 /OUT GND R
R3 Net-_D3-Pad1_ GND R
D3 Net-_D3-Pad1_ Net-_D3-Pad2_ LED
R4 Net-_D4-Pad1_ GND R
D4 Net-_D4-Pad1_ Net-_D4-Pad2_ LED
.end
